module zend

#include <php.h>
#include "v_bridge.h"
