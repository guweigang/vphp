module zend

pub const is_undef     = 0
pub const is_null      = 1
pub const is_false     = 2
pub const is_true      = 3
pub const is_long      = 4
pub const is_double    = 5
pub const is_string    = 6
pub const is_array     = 7
pub const is_object    = 8
